-0.8146782603592373,-0.9824024800333491,0.625340514212317,0.40790511960456777,0
0.9837290646229175,-0.37799078342032866,-0.05114904228682282,0.27449754699190976,0
-0.761488311113075,-0.9266300213533616,-0.7126869388914938,0.9834560407317621,0
-0.5581134912041716,0.14278019261775698,0.7463448113836775,0.2380178621716007,0
-0.5464100317311327,-0.7911795503814996,0.9589472112012545,0.6324435049805628,0
-0.08043054658606974,-0.27707093184759346,0.4075955630340333,-0.33852730792030017,0
-0.05254221026733097,-0.6663224259766034,0.41842864999347107,-0.62799737073745,0
0.24861154911019323,-0.23871792126876135,0.3498452217048582,-0.8474315947024642,0
-0.6528152499985183,0.3496795393519927,-0.05111280198117085,0.9895952669743842,0
-0.9395661714167138,0.9856894098072364,-0.44423226446396713,0.9661080729314995,0
0.5772993139080442,0.9903878442677012,-0.18994689963566813,-0.13370241425459528,0
0.7845128232324636,-0.6330688462097771,-0.71303914370847,0.17291896080719504,0
0.20295245773978454,0.38174240832579076,0.4769982770365404,0.44646922712235493,0
0.12023872042138639,-0.8407862370227088,0.2879206862637478,-0.4851751634835191,0
0.8239561937750601,0.5858885157305964,-0.18568589249337508,0.7598035485036725,0
0.9715488455458099,-0.9695464495543287,-0.10891893112509532,0.14872129311612214,0
0.732073395063354,-0.6022117736379007,-0.5839549468313681,0.37718640239916845,0
-0.1689152456400811,0.8321255362966962,-0.08693614715381481,0.8393222990030713,0
0.6602777239193249,0.24705765067446706,0.5083977283506007,-0.9410144993516523,0
-0.25207479454553705,-0.6748640851678367,0.4043772362289131,-0.036286192635294645,0
0.8759948526031347,0.0700176850813039,-0.722079856311082,0.04110473695188133,0
-0.2621113724282713,0.7409750669302422,-0.07638028634253846,0.7246296268810106,0
0.5277428098195764,0.37620036789357236,-0.48931974678785806,0.3618350594049087,0
-0.15535634797180942,-0.006140359162469133,0.23197239882314413,-0.150950468828565,0
-0.03148440020823351,-0.3874822929205717,0.00022104020579050143,0.5524905199922889,0
0.14052491674341971,-0.7919800612480123,-0.8632724832626355,0.16580197357208926,0
0.9729896655910957,0.0053302011801303895,0.9253127724794976,-0.6252576683914173,0
0.588372634197968,-0.8942363925315118,0.19660311904990757,-0.5126913223426706,0
-0.3785138124237495,0.10981764341118683,-0.12963773274731016,0.19850437276649124,0
-0.32682116764242886,-0.24050286297647383,-0.6736877340591882,0.3881763636468898,0
0.5868946449047345,0.34411643809039427,0.6635060779634316,0.43448293161251184,0
-0.4637329728618842,-0.5353894199221394,-0.7994632305427891,0.12857425312313042,0
0.9896436902244496,-0.4183351107701123,0.8484852708874924,-0.6511099835411929,0
0.5921651961950489,-0.8923801225845702,-0.5251445349470922,-0.18095403952236477,0
0.8731168676362269,0.7651164470943725,0.6434571273248411,0.590778663881449,0
-0.807482965926072,0.949461946806736,0.5178073539011352,0.08107090210826096,0
0.6181171029664363,-0.1853912069551853,0.4211917878622975,-0.9372030485888523,0
-0.7346826070967114,0.2799265697308535,0.7377563991587568,0.5119326429876883,0
-0.6110744430834458,-0.8097393831194213,-0.818779317519684,0.5361413636076202,0
0.7755892617373963,0.7400467735954719,0.5908744527729621,0.36863711336694127,0
-0.7072572592738573,-0.16341522471180037,-0.33018259237124714,0.604550585064261,0
-0.25848968120530946,-0.6102949646965601,0.5399389698156283,0.60794391609944,0
0.1179409422292832,0.4827872198616867,0.7158966637784692,0.9876825823126127,0
-0.16281738956090153,0.5957179338658816,0.5962390519454284,-0.7289544906391245,0
0.480943123328762,0.9428082934327262,0.2825431007442982,-0.7741325074615153,0
0.9464687548958308,-0.9722742578449561,0.5741576439775182,-0.7105528454796883,0
-0.8905134752037085,0.6841318608811886,0.8830781711387747,0.05332271533710631,0
0.3276797425909015,0.32142848827672754,-0.8432437442239193,0.912555615028086,0
0.5659362149906564,0.09569320780668877,-0.9536034508393092,0.29191450017078413,0
0.5142284047784598,0.2921352408338831,-0.6235253912860417,0.3941621320882007,0
0.5394498830743755,0.7244744467241109,-0.04694756656928356,0.050186044731995505,0
-0.8418383845726711,-0.2550730080358965,0.4382581086782613,0.9166688384292896,0
0.038171952940706744,0.7868559943399982,-0.10739995203959496,0.3083375838575344,0
0.0340873775815953,-0.9311131300028406,0.884428218088529,0.5854569484515715,0
-0.39280570053023856,-0.29388614982231664,0.07103831572633101,0.8446952090118001,0
-0.47534387601962624,0.4030324976068058,0.472650543239459,0.768591005410987,0
0.12759807342566964,-0.7263392720940518,-0.9793885112945453,-0.052630118663506975,0
0.00927762337950977,0.19093221056976972,0.5790576722383434,-0.05844065912256324,0
0.41157347102384634,-0.9866603216969736,0.2670622539581231,-0.06770755710021303,0
-0.04729462022737296,-0.8378950442046826,-0.9764229766848977,0.8828388861024188,0
0.2652990301868883,-0.09656422522320707,0.1741373081684623,0.07526617769283295,0
-0.6994648790379681,-0.311860342658542,0.8291293106692699,0.5824672952890213,0
0.7801361895077898,-0.8766955417240461,-0.05001125090081482,0.34917734733587946,0
0.4236914520694097,-0.5913650771425623,0.8487441138439742,-0.537570204228434,0
0.5557970943018451,0.22280753665666242,-0.7092903793752674,0.7929028537496805,0
0.6566846618759987,-0.34514923890132,-0.5720699990111642,0.08585018373629771,0
-0.2517977036491226,0.11635603658116422,-0.7674878525571653,0.9143798596474872,0
0.8107849520839274,0.9263668279752795,0.24496515870419788,-0.8668786276820237,0
0.5385166759632427,-0.12299143292460468,0.24206940511393582,-0.9514744745923243,0
0.0441855198491643,0.6672502800577589,-0.7608411246919788,0.13989887256545264,0
-0.23958315379161044,0.4740168393934665,0.39853410760202235,-0.8020013893558411,0
0.038171952940706744,0.7868559943399982,-0.05114904228682282,0.27449754699190976,0
-0.18322226500349645,0.5199135062426163,-0.8576330760886879,0.9876825823126127,0
-0.18322226500349645,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,0
-0.19076963390391882,0.5199135062426163,-0.8576330760886879,-0.36159484832566235,0
-0.18322226500349645,0.5199135062426163,-0.8576330760886879,0.9876825823126127,0
-0.18322226500349645,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,37
-0.19076963390391882,0.5199135062426163,-0.8576330760886879,-0.36159484832566235,38
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,46
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.052630118663506975,31
-0.18322226500349645,0.5907744041571028,-0.8576330760886879,0.768591005410987,0
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,34
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,33
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.052630118663506975,37
-0.19076963390391882,0.5957179338658816,0.5962390519454284,-0.7289544906391245,0
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.33793179963228814,40
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.052630118663506975,41
-0.18322226500349645,0.5907744041571028,-0.8576330760886879,-0.05035247491201984,36
-0.19269911704030884,0.5213579012823353,-0.8576330760886879,-0.5126913223426706,37
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,39
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,40
-0.18322226500349645,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,50
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.052630118663506975,21
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,38
-0.18322226500349645,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,45
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,0.40790511960456777,0
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.052630118663506975,41
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.36159484832566235,40
-0.18322226500349645,0.5907744041571028,-0.8576330760886879,0.3881763636468898,0
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.052630118663506975,28
-0.18322226500349645,0.5907744041571028,0.5741576439775182,-0.7105528454796883,0
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.052630118663506975,37
-0.19076963390391882,0.5907744041571028,-0.8576330760886879,-0.052630118663506975,31
