11
-0.6242355062709293,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,51
-0.2548597909717818,0.6732527641816939,-0.8975174536762058,-0.31478386254215707,75
-0.2548597909717818,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,70
-0.2548597909717818,0.8675694905501019,-0.5435142648368467,-0.06021783134623249,50
-0.2548597909717818,0.8675694905501019,-1.0745654464705994,-0.31478386254215707,63
-0.2548597909717818,0.6732527641816939,-0.8458665536291754,-0.31478386254215707,68
-0.2548597909717818,0.8675694905501019,-0.8975174536762058,-0.31478386254215707,60
-0.2548597909717818,0.8675694905501019,-0.5435142648368467,-0.31478386254215707,70
-0.2548597909717818,0.8675694905501019,-0.5435142648368467,-0.31478386254215707,66
-0.2548597909717818,1.125884076372659,-0.8975174536762058,-0.31478386254215707,76
-0.2548597909717818,0.8675694905501019,-0.8975174536762058,-0.2936471948015749,77
-0.2548597909717818,0.8675694905501019,-0.5435142648368467,-0.31478386254215707,72
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.31478386254215707,74
-0.2548597909717818,0.877514103976044,-0.6688043868506017,-0.31478386254215707,63
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.31478386254215707,69
-0.2548597909717818,0.8675694905501019,-0.5435142648368467,-0.06021783134623249,75
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.31478386254215707,74
-0.2548597909717818,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,68
-0.2548597909717818,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,72
-0.2548597909717818,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,71
-0.2548597909717818,1.125884076372659,-0.8975174536762058,-0.31478386254215707,70
-0.2548597909717818,0.8675694905501019,-0.5435142648368467,-0.31478386254215707,67
-0.2548597909717818,0.8675694905501019,-0.5266337414513725,-0.4064282184720165,59
-0.2548597909717818,0.8675694905501019,-0.8975174536762058,-0.31478386254215707,74
-0.2548597909717818,0.8675694905501019,-0.8975174536762058,-0.31478386254215707,74
-0.6242355062709293,1.125884076372659,-0.8649689913693525,-0.31478386254215707,68
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.31478386254215707,72
-0.2548597909717818,0.8675694905501019,-0.5435142648368467,-0.06021783134623249,74
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.31478386254215707,63
-0.2548597909717818,0.8675694905501019,-0.8168910066990992,-0.31478386254215707,63
-0.2548597909717818,0.6732527641816939,-0.6688043868506017,-0.31478386254215707,63
-0.6242355062709293,1.125884076372659,-0.4090467039036283,-0.06021783134623249,63
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.48680738412331825,63
-0.6242355062709293,0.6732527641816939,-0.6688043868506017,-0.4064282184720165,63
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.618464685441283,63
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.4064282184720165,63
-0.2548597909717818,0.6053465813871026,-0.5435142648368467,-0.06021783134623249,63
-0.30883291749164304,1.125884076372659,-0.8458665536291754,-0.48680738412331825,64
-0.6242355062709293,1.125884076372659,-0.3438235898527883,-0.31478386254215707,64
-0.2548597909717818,0.8675694905501019,-0.4090467039036283,-0.31478386254215707,64
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.48680738412331825,64
-0.2548597909717818,0.6732527641816939,-0.8458665536291754,-0.2991132043883876,64
-0.6242355062709293,1.125884076372659,-0.8458665536291754,-0.48680738412331825,64
-0.6242355062709293,1.125884076372659,-0.8458665536291754,-0.06021783134623249,64
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.31478386254215707,65
-0.6242355062709293,1.125884076372659,-0.6688043868506017,-0.48680738412331825,65
-0.2548597909717818,0.6732527641816939,-0.8458665536291754,-0.31478386254215707,65
-0.6242355062709293,0.6732527641816939,-0.6688043868506017,-0.4064282184720165,65
-0.2548597909717818,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,65
-0.6242355062709293,1.125884076372659,-0.6688043868506017,-0.48680738412331825,65
-0.11796767456636381,0.8675694905501019,-0.6688043868506017,-0.48680738412331825,65
-0.2548597909717818,0.8675694905501019,-0.8975174536762058,-0.31478386254215707,66
-0.2548597909717818,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,66
-0.2548597909717818,0.6732527641816939,-0.6688043868506017,-0.4064282184720165,66
-0.6242355062709293,0.6053465813871026,-0.8975174536762058,-0.31478386254215707,66
-0.2548597909717818,0.6732527641816939,-0.8458665536291754,-0.48680738412331825,66
-0.6242355062709293,0.6732527641816939,-0.8458665536291754,-0.48680738412331825,66
-0.2548597909717818,0.8675694905501019,-0.6688043868506017,-0.03082578600969356,67
-0.6242355062709293,1.125884076372659,-0.8458665536291754,-0.31478386254215707,67
-0.6734206646825089,1.125884076372659,-0.8458665536291754,-0.31478386254215707,67
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.31478386254215707,67
-0.30883291749164304,0.6053465813871026,-0.8975174536762058,-0.31478386254215707,67
-0.6242355062709293,1.125884076372659,-0.8458665536291754,-0.4064282184720165,67
-0.11796767456636381,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,67
-0.2548597909717818,0.6732527641816939,-0.6688043868506017,-0.4064282184720165,67
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.31478386254215707,68
-0.30883291749164304,0.6053465813871026,-0.8975174536762058,-0.31478386254215707,68
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.31478386254215707,68
-0.2548597909717818,0.6053465813871026,-0.8975174536762058,-0.31478386254215707,68
-0.2548597909717818,0.6732527641816939,-0.8458665536291754,-0.48680738412331825,68
-0.2548597909717818,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,69
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.31478386254215707,69
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.31478386254215707,69
-0.6242355062709293,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,69
-0.6242355062709293,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,69
-0.2548597909717818,0.6732527641816939,-0.6688043868506017,-0.4064282184720165,69
-0.6242355062709293,1.125884076372659,-0.6688043868506017,-0.31478386254215707,69
-0.30883291749164304,0.6053465813871026,-0.8975174536762058,-0.4064282184720165,69
-0.6242355062709293,1.125884076372659,-0.8458665536291754,-0.618464685441283,69
-0.2548597909717818,0.8675694905501019,-0.4090467039036283,-0.31478386254215707,69
-0.2548597909717818,0.877514103976044,-0.6688043868506017,-0.31478386254215707,70
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.31478386254215707,70
-0.2548597909717818,0.6053465813871026,-0.5435142648368467,-0.06021783134623249,70
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.31478386254215707,70
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.31478386254215707,71
-0.6242355062709293,1.125884076372659,-0.8458665536291754,-0.48680738412331825,72
-0.2548597909717818,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,73
-0.6242355062709293,1.125884076372659,-0.8975174536762058,-0.31478386254215707,73
-0.2548597909717818,0.8675694905501019,-0.8975174536762058,-0.2991132043883876,73
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.31478386254215707,73
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.4064282184720165,73
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.48680738412331825,73
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.4064282184720165,74
-0.2548597909717818,0.6732527641816939,-0.8458665536291754,-0.31478386254215707,74
-0.2548597909717818,0.8675694905501019,-0.5435142648368467,-0.06021783134623249,74
-0.2548597909717818,0.8675694905501019,-0.6688043868506017,-0.31478386254215707,74
-0.2548597909717818,0.8675694905501019,-0.8975174536762058,-0.31478386254215707,75
-0.2548597909717818,0.6732527641816939,-0.8458665536291754,-0.2991132043883876,76
-0.2548597909717818,0.8675694905501019,-0.8458665536291754,-0.31478386254215707,77
-0.2548597909717818,0.8675694905501019,-0.8975174536762058,-0.31478386254215707,77
